// $Id: $
// File name:   test.sv
// Created:     4/18/2016
// Author:      Pradeep Kumar Lam
// Lab Section: 337-03
// Version:     1.0  Initial Design Entry
// Description: This is for testing ideas/concepts.



