// $Id: $
// File name:   writeController.sv
// Created:     4/24/2016
// Author:      Pradeep Kumar Lam
// Lab Section: 337-03
// Version:     1.0  Initial Design Entry
// Description: This is what controls the writing of data to the fpga.
